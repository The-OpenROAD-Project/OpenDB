#################################################################################
#										#
# 	Version		:	5.5						#
# 	Last updated 	:	04/05/99					#
#										#
#################################################################################

VERSION 5.5 ;
NAMESCASESENSITIVE ON ;
NOWIREEXTENSIONATPIN ON ;
BUSBITCHARS "<>" ;
DIVIDERCHAR ":" ;
MANUFACTURINGGRID 3.5 ;
USEMINSPACING OBS OFF ;
USEMINSPACING PIN ON ;
CLEARANCEMEASURE EUCLIDEAN ;
CLEARANCEMEASURE MAXXY ;

UNITS
  TIME NANOSECONDS 100 ;
  CAPACITANCE PICOFARADS 10 ;
  RESISTANCE OHMS 10000 ;
  POWER MILLIWATTS 10000 ;
  CURRENT MILLIAMPS 10000 ;
  VOLTAGE VOLTS 1000 ;
  DATABASE MICRONS 1000 ;
  FREQUENCY MEGAHERTZ 10 ;
END UNITS

PROPERTYDEFINITIONS
	LIBRARY NAME STRING "Cadence96" ;
	LIBRARY intNum  INTEGER 20 ;
	LIBRARY realNum REAL 21.22 ;
	LAYER lsp STRING ;
	LAYER lip INTEGER ;
	LAYER lrp REAL ;
	VIA stringProperty STRING ;
	VIA realProperty REAL ;
	VIA COUNT INTEGER RANGE 1 100 ;
	VIARULE vrsp STRING ;
	VIARULE vrip INTEGER ;
	VIARULE vrrp REAL ;
	NONDEFAULTRULE ndrsp STRING ;
	NONDEFAULTRULE ndrip INTEGER ;
	NONDEFAULTRULE ndrrp REAL ;
	MACRO stringProp STRING ;
	MACRO integerProp INTEGER ;
	MACRO WEIGHT REAL RANGE 1.0 100.0 ;
	PIN TYPE STRING ;
	PIN intProp INTEGER ;
	PIN realProp REAL ;
END PROPERTYDEFINITIONS

LAYER POLYS
	TYPE MASTERSLICE ;
	PROPERTY lsp "top" lip 1 lrp 2.3 ;
END POLYS

LAYER CUT01
	TYPE CUT ;
        SPACING 0.35 ADJACENTCUTS 3 WITHIN 0.25 ;
	PROPERTY lip 5 ;
END CUT01

LAYER RX
	TYPE ROUTING ;
	PITCH 1.8 ;
	OFFSET 0.9 ;
	WIDTH 1 ;
        AREA 34.1 ;
        MINIMUMCUT 2 WIDTH 2.5 ;
	SPACING 0.6 ;
	SPACING 0.18 LENGTHTHRESHOLD 0.9 ;
	SPACING 0.4 RANGE 0.1 0.12 ;
	SPACING 0.32 RANGE 1.01 2000.0 USELENGTHTHRESHOLD ;
        SPACING 0.1 RANGE 0.1 0.1 INFLUENCE 2.01 RANGE 2.1 10000.0 ;
        SPACING 0.44 RANGE 1.0 1.0 INFLUENCE 1.01 ;
	SPACING 0.33 RANGE 1.01 20.0 INFLUENCE 1.01 ;
	SPACING 0.7 RANGE 0.3 0.15 USELENGTHTHRESHOLD ;
	SPACING 0.5 ;
	SPACING 0.6 RANGE 4.5 6.12 RANGE 3.0 3.1 ;
        SPACING 4.3 RANGE 0.1 0.1 INFLUENCE 3.81 RANGE 0.1 0.2 ;
        SPACING 0.53 LENGTHTHRESHOLD 0.45 RANGE 0 0.1 ;
	DIRECTION HORIZONTAL ;
	WIREEXTENSION 0.75 ;
	RESISTANCE RPERSQ 0.103 ;
	CAPACITANCE CPERSQDIST 0.000156 ;
	HEIGHT 9 ;
	THICKNESS 1 ;
	SHRINKAGE 0.1 ;
        SLOTWIREWIDTH 5 ;
        SLOTWIRELENGTH 4 ;
        SLOTWIDTH 6 ;
        SLOTLENGTH 5 ;
        MAXADJACENTSLOTSPACING 45 ;
        MAXCOAXIALSLOTSPACING 55 ;
        SPLITWIREWIDTH 5 ;
        MINIMUMDENSITY 4 ;
        MAXIMUMDENSITY 10 ;
#        DENSITYCHECKWINDOW 4 5 ;
        DENSITYCHECKSTEP 2 ;
        FILLACTIVESPACING 4 ;
	CAPMULTIPLIER 1 ;
	EDGECAPACITANCE 0.00005 ;
        ANTENNAMODEL OXIDE1 ;
	ANTENNAAREAFACTOR 1 ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAAREARATIO 4.6 ;
        ANTENNAAREARATIO 7.6 ;
        ANTENNADIFFAREARATIO 4.7 ;
        ANTENNADIFFAREARATIO PWL ( ( 5.4 5.4 ) ( 6.5 6.5 ) ( 7.5 7.5 ) ) ;
        ANTENNACUMAREARATIO 6.7 ;
        ANTENNACUMDIFFAREARATIO 4.5 ;
        ANTENNACUMDIFFAREARATIO PWL ( ( 5.4 5.4 ) ( 6.5 6.5 ) ( 7.5 7.5 ) ) ;
        ANTENNAAREAFACTOR 6.5 ;
        ANTENNAAREAFACTOR 6.5 DIFFUSEONLY ;
        ANTENNASIDEAREARATIO 6.5 ;
        ANTENNADIFFSIDEAREARATIO 6.5 ;
        ANTENNADIFFSIDEAREARATIO PWL ( ( 5.4 5.4 ) ( 6.5 6.5 ) ( 7.5 7.5 ) ) ;
        ANTENNACUMSIDEAREARATIO 4.5 ;
        ANTENNACUMSIDEAREARATIO 7.5 ;
        ANTENNACUMDIFFSIDEAREARATIO 4.6 ; 
        ANTENNACUMDIFFSIDEAREARATIO PWL ( ( 5.4 5.4 ) ( 6.5 6.5 ) ( 7.5 7.5 ) ) ;
        ANTENNASIDEAREAFACTOR 6.5 ;
        ANTENNASIDEAREAFACTOR 7.5 DIFFUSEONLY ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAMODEL OXIDE4 ;
	PROPERTY lsp "rxlay" lip 3 lrp 1.2 ;
        CURRENTDEN 1E3 ;
#        CURRENTDEN ( 1E3 4E5 ) ;
	ACCURRENTDENSITY PEAK
	  FREQUENCY 1E6 100E6 ;
	  TABLEENTRIES 0.5E-6 0.4E-6 ;
	ACCURRENTDENSITY AVERAGE 5.5 ;
	ACCURRENTDENSITY RMS
	  FREQUENCY 100E6 400E6 800E6 ;
	  WIDTH     0.4 0.8 10.0 50.0 100.0 ;
	  TABLEENTRIES
	    2.0E-6 1.9E-6 1.8E-6 1.7E-6 1.5E-6
	    1.4E-6 1.3E-6 1.2E-6 1.1E-6 1.0E-6
	    0.9E-6 0.8E-6 0.7E-6 0.6E-6 0.4E-6 ;
	DCCURRENTDENSITY AVERAGE
	  WIDTH 20.0 50.0 ;
	  TABLEENTRIES 0.6E-6 0.5E-6 ;
END RX

LAYER CUT12
	TYPE CUT ;
	SPACING 0.7 LAYER RX ;
        SPACING 0.22 ADJACENTCUTS 4 WITHIN 0.25 ;
        # 5.4
        ANTENNAMODEL OXIDE1 ;
        ANTENNAMODEL OXIDE2 ;
        ANTENNAMODEL OXIDE3 ;
        ANTENNAMODEL OXIDE4 ;
        ANTENNAAREAFACTOR 5.4 ;
        ANTENNADIFFAREARATIO 6.5 ;
        ANTENNADIFFAREARATIO PWL ( ( 5.4 5.4 ) ( 6.5 6.5 ) ( 7.5 7.5 ) ) ;
        ANTENNACUMDIFFAREARATIO PWL ( ( 5.4 5.4 ) ( 6.5 6.5 ) ( 7.5 7.5 ) ) ;
        ANTENNACUMDIFFAREARATIO 5.6 ;
        ANTENNAAREARATIO 5.6 ;
        ANTENNACUMAREARATIO 6.7 ;
	ACCURRENTDENSITY PEAK
	  FREQUENCY 1E6 100E6 ;
	  TABLEENTRIES 0.5E-6 0.4E-6 ;
	ACCURRENTDENSITY AVERAGE 5.5 ;
	ACCURRENTDENSITY RMS
	  FREQUENCY 100E6 400E6 800E6 ;
	  WIDTH     0.4 0.8 10.0 50.0 100.0 ;
	  TABLEENTRIES
	    2.0E-6 1.9E-6 1.8E-6 1.7E-6 1.5E-6
	    1.4E-6 1.3E-6 1.2E-6 1.1E-6 1.0E-6
	    0.9E-6 0.8E-6 0.7E-6 0.6E-6 0.4E-6 ;
	DCCURRENTDENSITY AVERAGE
          CUTAREA 2.0 5.0 ; 
          TABLEENTRIES 0.5E-6 0.4E-6 ;
	DCCURRENTDENSITY AVERAGE 4.9 ;
END CUT12

LAYER PC
	TYPE ROUTING ;
	WIDTH 1 ;
	WIREEXTENSION 0.4 ; #should be ignored
	PITCH 1.8 ;
	SPACING 0.6 ;
	DIRECTION VERTICAL ;
	RESISTANCE RPERSQ PWL ( ( 1 0.103 ) ( 10 4.7 ) ) ;
	CAPACITANCE CPERSQDIST PWL ( ( 1 0.000156 ) ( 10 0.001 ) ) ;
        ANTENNAAREARATIO 5.4 ;
        ANTENNADIFFAREARATIO 6.5 ;
        ANTENNACUMAREARATIO 7.5 ;
        ANTENNACUMDIFFAREARATIO PWL ( ( 5.0 5.1 ) ( 6.0 6.1 ) ) ;
        ANTENNAAREAFACTOR 4.5 ;
        ANTENNASIDEAREARATIO 6.5 ;
        ANTENNADIFFSIDEAREARATIO PWL ( ( 7.0 7.1 ) ( 7.2 7.3 ) ) ;  
        ANTENNACUMSIDEAREARATIO 7.4 ;
        ANTENNACUMDIFFSIDEAREARATIO PWL ( ( 8.0 8.1 ) ( 8.2 8.3 ) ( 8.4 8.5 )
             ( 8.6 8.7 ) ) ;
        ANTENNASIDEAREAFACTOR 9.0 DIFFUSEONLY ;

        ACCURRENTDENSITY PEAK
          FREQUENCY 1E6 100E6 ;
          CUTAREA 5.6 8.5 8.1 4.5 ;
          TABLEENTRIES 0.5E-6 0.4E-6 ;
	DCCURRENTDENSITY AVERAGE
	  WIDTH 20.0 50.0 100.0 ;
	  TABLEENTRIES 1.0E-6 0.7E-6 0.5E-6 ;
END PC

LAYER CA
	TYPE CUT ;
	DCCURRENTDENSITY AVERAGE
	  CUTAREA   2.0 5.0 10.0 ;
	  TABLEENTRIES 0.6E-6 0.5E-6 0.4E-6 ; 
END CA

LAYER M1
	TYPE ROUTING ;
	WIDTH 1 ;
	WIREEXTENSION 7 ;
	PITCH 1.8 ;
	DIRECTION HORIZONTAL ;
	RESISTANCE RPERSQ 0.103 ;
	CAPACITANCE CPERSQDIST 0.000156 ;
        ANTENNACUMAREARATIO 300 ;
        ANTENNACUMDIFFAREARATIO 600 ;
        SPACINGTABLE
          PARALLELRUNLENGTH 0.00 0.50 3.00 5.00
            WIDTH 0.00      0.15 0.15 0.15 0.15
            WIDTH 0.25      0.15 0.20 0.20 0.20
            WIDTH 1.50      0.15 0.50 0.50 0.50
            WIDTH 3.00      0.15 0.50 1.00 1.00
            WIDTH 5.00      0.15 0.50 1.00 2.00 ;
        SPACINGTABLE
          INFLUENCE
            WIDTH 1.5 WITHIN 0.5 SPACING 0.5
            WIDTH 3.0 WITHIN 1.0 SPACING 1.0
            WIDTH 5.0 WITHIN 2.0 SPACING 2.0 ;
        ACCURRENTDENSITY AVERAGE 5.5 ;
        DCCURRENTDENSITY AVERAGE 4.9 ;
END M1

LAYER V1
	TYPE CUT ;
	SPACING 0.6 LAYER CA ;
END V1

LAYER M2
	TYPE ROUTING ;
	WIDTH 0.9 ;
	WIREEXTENSION 8 ;
	PITCH 1.8 ;
	SPACING 0.9 ;
        SPACING 0.28 ;
        SPACING 0.24 LENGTHTHRESHOLD 1.0 ;
        SPACING 0.32 RANGE 1.01 9.99 USELENGTHTHRESHOLD ;
        SPACING 0.5 RANGE 10.0 1000.0 ;
        SPACING 0.5 RANGE 10.0 1000.0 INFLUENCE 1.00 ;
        SPACING 0.5 RANGE 10.0 1000.0 INFLUENCE 1.0 RANGE .28 1.0 ;
        SPACING 0.5 RANGE 3.01 4.0 RANGE 4.01 5.0 ;
        SPACING 0.4 RANGE 3.01 4.0 RANGE 5.01 1000.0 ;
	DIRECTION VERTICAL ;
	RESISTANCE RPERSQ 0.0608 ;
	CAPACITANCE CPERSQDIST 0.000184 ;
END M2

LAYER V2
	TYPE CUT ;
END V2

LAYER M3
	TYPE ROUTING ;
	WIDTH 0.9 ;
	WIREEXTENSION 8 ;
	PITCH 1.8 ;
	SPACING 0.9 ;
	DIRECTION HORIZONTAL ;
	RESISTANCE RPERSQ 0.0608 ;
	CAPACITANCE CPERSQDIST 0.000184 ;
END M3

LAYER M4
        TYPE ROUTING ;
        PITCH 5.4 ;
        WIDTH 5.4 ;
        DIRECTION VERTICAL ;
        DIRECTION HORIZONTAL ;
        # 2 via cuts required for m4 > 0.50 um when connecting from m3
        MINIMUMCUT 2 WIDTH 0.50 ;
        # 2 via cuts required for m4 > 0.70 um when connecting from m5
        MINIMUMCUT 2 WIDTH 0.70 FROMBELOW ;
        # 4 via cuts are required for m4 > 1.0 um when connecting from m3 or m5
        MINIMUMCUT 4 WIDTH 1.0 FROMABOVE ;
        # 2 via cuts are required if m4 > 1.1 um wide and m4 > 20.0 um long,
        # and the via cut is < 5.0 um away from the wide wire
        MINIMUMCUT 2 WIDTH 1.1 LENGTH 20.0 WITHIN 5.0 ;
        MINIMUMCUT 2 WIDTH 1.1 FROMABOVE LENGTH 20.0 WITHIN 5.0 ;
        MINENCLOSEDAREA 0.30 ; # donut hole must be >= 0.30 um^2
        MINENCLOSEDAREA 0.40 WIDTH 0.15 ; # hole area >= 0.40 um^2 when w<=0.15
        MINENCLOSEDAREA 0.80 WIDTH 0.50 ; # hole area >= 0.80 um^2 when w<=0.55
        MAXWIDTH 10.0 ;
        MINWIDTH 0.15 ;
        PROTRUSIONWIDTH 0.30 LENGTH 0.60 WIDTH 1.20 ;
        MINSTEP .20 ;
END M4

LAYER M5
        TYPE ROUTING ;
        PITCH 5.4 ;
        WIDTH 4.0 ;
        DIRECTION VERTICAL ;
        MINIMUMCUT 2 WIDTH 0.70 ;
        MINIMUMCUT 4 WIDTH 1.0 FROMABOVE ;
        MINIMUMCUT 2 WIDTH 1.1 LENGTH 20.0 WITHIN 5.0 ;
        MINIMUMCUT 5 WIDTH 0.5  ;
END M5

LAYER implant1
        TYPE IMPLANT ;
        WIDTH 0.50 ;
        SPACING 0.50 ;
        PROPERTY lrp 5.4 ;
END implant1
        
LAYER implant2
        TYPE IMPLANT ;
        WIDTH 0.50 ;
        SPACING 0.50 ;
        PROPERTY lsp "bottom" ;
END implant2

LAYER V3
	TYPE CUT ;
END V3

LAYER MT
	TYPE ROUTING ;
	WIDTH 0.9 ;
	PITCH 1.8 ;
	SPACING 0.9 ;
	DIRECTION VERTICAL ;
	RESISTANCE RPERSQ 0.0608 ;
	CAPACITANCE CPERSQDIST 0.000184 ;
END MT

layer OVERLAP
	TYPE OVERLAP ;
        PROPERTY lip 5 lsp "top" ;
        PROPERTY lrp 5.5 lsp "bottom" ;
END OVERLAP

MAXVIASTACK 4 RANGE m1 m7 ;

#layer VIRTUAL
#	TYPE OVIRTUAL ;
#END VIRTUAL

VIA IN1X
	TOPOFSTACKONLY 
	FOREIGN IN1X ;
	RESISTANCE 2 ;
	LAYER RX ;
	  RECT -0.7 -0.7 0.7 0.7 ;
	LAYER CUT12 ;
	  RECT -0.25 -0.25 0.25 0.25 ;
	LAYER PC ;
	  RECT -0.6 -0.6 0.6 0.6 ;
	PROPERTY stringProperty "DEFAULT" realProperty 32.33 COUNT 34 ;
END IN1X

VIA M1_M2 DEFAULT
	RESISTANCE 1.5 ;
	LAYER M1 ;
	  RECT -0.6 -0.6 0.6 0.6 ;
	LAYER V1 ;
	  RECT -0.45 -0.45 0.45 0.45 ;
	LAYER M2 ;
	  RECT -0.45 -0.45 0.45 0.45 ;
END M1_M2

VIA M2_M3 DEFAULT
	RESISTANCE 1.5 ;
	LAYER M2 ;
	  RECT -0.45 -0.9 0.45 0.9 ;
	LAYER V2 ;
	  RECT -0.45 -0.45 0.45 0.45 ;
	LAYER M3 ;
	  RECT -0.45 -0.45 0.45 0.45 ;
END M2_M3

VIA M2_M3_PWR 
	RESISTANCE 0.4 ;
	LAYER M2 ;
	  RECT -1.35 -1.35 1.35 1.35 ;
	LAYER V2 ;
	  RECT -1.35 -1.35 -0.45 1.35 ;
	  RECT 0.45 -1.35 1.35 -0.45 ;
	  RECT 0.45 0.45 1.35 1.35 ;
	LAYER M3 ;
	  RECT -1.35 -1.35 1.35 1.35 ;
END M2_M3_PWR

VIA M3_MT DEFAULT
	RESISTANCE 1.5 ;
	LAYER M3 ;
	  RECT -0.9 -0.45 0.9 0.45 ;
	LAYER V3 ;
	  RECT -0.45 -0.45 0.45 0.45 ;
	LAYER MT ;
	  RECT -0.45 -0.45 0.45 0.45 ;
END M3_MT

VIA VIACENTER12
  LAYER M1 ;
      RECT -4.6 -2.2 4.6 2.2 ;
  LAYER V1 ;
      RECT -3.1 -0.8 -1.9 0.8 ;
      RECT 1.9 -0.8 3.1 0.8 ;
  LAYER M2 ;
      RECT -4.4 -2.0 4.4 2.0 ;
  RESISTANCE 0.24 ; 
END VIACENTER12

VIA M2_TURN 
  LAYER M2 ;
      RECT -0.45 -0.45 0.45 0.45 ;
      RECT -4.4 -2.0 4.4 2.0 ;
END M2_TURN

VIARULE VIALIST12
  LAYER M1 ;
      DIRECTION VERTICAL ;
      OVERHANG 4.5 ;
      WIDTH 9.0 TO 9.6 ;
      METALOVERHANG 0.4 ;
  LAYER M2 ;
      DIRECTION HORIZONTAL ;
      WIDTH 3.0 TO 3.0 ;
      METALOVERHANG 0.3 ;
  VIA VIACENTER12 ;
  PROPERTY vrsp "new" vrip 1 vrrp 4.5 ;
END VIALIST12

VIARULE VIALIST1
  LAYER M1 ;
      DIRECTION VERTICAL ;
      WIDTH 9.0 TO 9.6 ;
      OVERHANG 4.5 ;
      METALOVERHANG 0.5 ;
  LAYER M1 ;
      DIRECTION HORIZONTAL ;
      WIDTH 3.0 TO 3.0 ;
      OVERHANG 5.5 ;
      METALOVERHANG 0.6 ;
  VIA VIACENTER12 ;
END VIALIST1
 

VIARULE VIAGEN12 GENERATE 
   LAYER M1 ;
	DIRECTION VERTICAL ;
	WIDTH 0.1 TO 19 ;
	OVERHANG 1.4 ;
	METALOVERHANG 1.0 ;
   LAYER M2 ;
	DIRECTION HORIZONTAL ;
	OVERHANG 1.4 ;
	METALOVERHANG 1.0 ;
        WIDTH 0.2 TO 1.9 ;
  LAYER M3 ;
      RECT -0.3 -0.3 0.3 0.3 ;
      SPACING 5.6 BY 7.0 ;
      RESISTANCE 0.5 ; 
  PROPERTY vrsp "new" vrip 1 vrrp 5.5 ;
END VIAGEN12

VIARULE VIAGEN1 GENERATE 
   LAYER M1 ;
	DIRECTION HORIZONTAL ;
	OVERHANG 1.4 ;
	METALOVERHANG 1.1 ;
	WIDTH 0.1 TO 1.9 ;
   LAYER M1 ;
	DIRECTION VERTICAL ;
	OVERHANG 1.5 ;
	METALOVERHANG 1.5 ;
        WIDTH 0.2 TO 2.9 ;
   LAYER M1 ;
        RECT ( 1 1 ) ( 1 1 ) ;
        SPACING 0.3 BY 4.5 ;
  PROPERTY vrsp "new" vrip 1 vrrp 5.5 ;
END VIAGEN1

VIARULE via12 GENERATE
  LAYER m1 ;
        ENCLOSURE 0.05 0.005 ; # 2 sides need >= 0.05, 2 other sides >= 0.005
        WIDTH 1.0 TO 100.0 ;   # for m1 between 1 to 100 um wide
  LAYER m2 ;
        ENCLOSURE 0.05 0.005 ; # 2 sides need >= 0.05, 2 other sides >= 0.005
        WIDTH 1.0 TO 100.0 ;   # for m1 between 1 to 100 um wide
  LAYER cut12 ;
        RECT -0.07 -0.07 0.07 0.07 ; # cut is .14 by .14
        SPACING 0.16 BY 0.16 ;
END via12


NONDEFAULTRULE RULE1
    LAYER RX
	WIDTH 10.0 ;
	SPACING 2.2 ;
	WIREEXTENSION 6 ;
        RESISTANCE RPERSQ 6.5 ;
        CAPACITANCE CPERSQDIST 6.5 ;
        EDGECAPACITANCE 6.5 ;
    END RX
    LAYER PC
	WIDTH 10.0 ;
	SPACING 2.2 ;
        CAPACITANCE CPERSQDIST 6.5 ;
    END PC

    LAYER M1
        WIDTH 10.0 ;
	SPACING 2.2 ;
        RESISTANCE RPERSQ 6.5 ;
    END M1
     
    VIA nd1VIARX0
         DEFAULT
         TOPOFSTACKONLY
	 FOREIGN IN1X ;
	 RESISTANCE 0.2 ;
         PROPERTY realProperty 2.3 ;
	 LAYER RX ;
	  RECT -3 -3 3 3 ;
	 LAYER CUT12 ;
	  RECT -1.0 -1.0 1.0 1.0 ;
	 LAYER PC ;
	  RECT -3 -3 3 3 ;
    END nd1VIARX0

    VIA nd1VIA01
        FOREIGN IN1X 5.6 5.3 E ;
	RESISTANCE 0.2 ;
	LAYER PC ;
	  RECT -3 -3 3 3 ;
          RECT -5 -5 5 5 ;
	LAYER CA ;
	  RECT -1.0 -1.0 1.0 1.0 ;
	LAYER M1 ;
	  RECT -3 -3 3 3 ;
    END nd1VIA01
    VIA nd1VIA12

	 RESISTANCE 0.2 ;
	 LAYER M1 ;
	  RECT -3 -3 3 3 ;
	 LAYER V1 ;
          RECT -1.0 -1.0 1.0 1.0 ;
         LAYER M2 ;
	  RECT -3 -3 3 3 ;
     END nd1VIA12
				    
     SPACING
	 SAMENET
	  CUT01 RX 0.1 STACK ;
     END SPACING
     PROPERTY ndrsp "single" ndrip 1 ndrrp 6.7 ;
END RULE1

UNIVERSALNOISEMARGIN 0.1 20 ;
EDGERATETHRESHOLD1 0.1 ;
EDGERATETHRESHOLD2 0.9 ;
EDGERATESCALEFACTOR 1.0 ;

NOISETABLE 1 ;
	EDGERATE 20 ;
	OUTPUTRESISTANCE 3 ;
	VICTIMLENGTH 25 ;
	VICTIMNOISE 10 ;
#        CORRECTIONFACTOR 3 ;
#        OUTPUTRESISTANCE 5 ;
END NOISETABLE

#CORRECTIONTABLE 1 ;
#	EDGERATE 20 ;
#	OUTPUTRESISTANCE 3 ;
#	VICTIMLENGTH 25 ;
#	CORRECTIONFACTOR 10.5 ;
#        OUTPUTRESISTANCE 5.4 ;
#END CORRECTIONTABLE

SPACING
	SAMENET CUT01 CA 1.5 ;
	SAMENET CA V1 1.5 STACK ;
	SAMENET M1 M1 3.5 STACK ;
	SAMENET V1 V2 1.5 STACK ;
	SAMENET M2 M2 3.5 STACK ;
	SAMENET V2 V3 1.5 STACK ;
END SPACING

MINFEATURE 0.1 0.1 ;

DIELECTRIC 0.000345 ;

IRDROP 
	TABLE DRESHI
		0.0001 -0.7 0.001 -0.8 0.01 -0.9 0.1 -1.0 ;
	TABLE DRESLO
		0.0001 -1.7 0.001 -1.6 0.01 -1.5 0.1 -1.3 ;
	TABLE DNORESHI
		0.0001 -0.6 0.001 -0.7 0.01 -0.9 0.1 -1.1 ;
	TABLE DNORESLO
		0.0001 -1.5 0.001 -1.5 0.01 -1.4 0.1 -1.4 ;
END IRDROP

SITE  COVER
        CLASS PAD ;
        SYMMETRY R90 ;
        SIZE 10.000 BY 10.000 ;
END  COVER

SITE  IO
        CLASS PAD ;
        SIZE 80.000 BY 560.000 ;
END  IO

SITE  CORE
        CLASS CORE ;
        SIZE 0.700 BY 8.400 ;
END  CORE

SITE CORE1
  	CLASS CORE ;
    	SYMMETRY X ;
      	SIZE 67.2 BY 6 ;
END CORE1

SITE MRCORE
#	CLASS VIRTUAL ;
	CLASS CORE ;
	SIZE 3.6 BY 28.8 ;
	SYMMETRY  Y  ;
END MRCORE

SITE IOWIRED
	CLASS PAD ;
	SIZE 57.6 BY 432 ;
END IOWIRED

SITE IMAGE
	CLASS CORE ;
	SIZE 1 BY 1 ;
END IMAGE

ARRAY M7E4XXX
    SITE CORE            -5021.450 -4998.000 N DO 14346 BY 595 STEP 0.700 16.800 ;
    SITE CORE            -5021.450 -4989.600 FS DO 14346 BY 595 STEP 0.700 16.800 ;
    SITE IO              6148.800 5800.000 E DO 1 BY 1 STEP 0.000 0.000 ;
    SITE IO              6148.800 3240.000 E DO 1 BY 1 STEP 0.000 0.000 ;
    SITE COVER           -7315.000 -7315.000 N DO 1 BY 1 STEP 0.000 0.000 ;
    SITE COVER           7305.000 7305.000 N DO 1 BY 1 STEP 0.000 0.000 ;
    CANPLACE COVER           -7315.000 -7315.000 N DO 1 BY 1 STEP 0.000 0.000 ;
    CANPLACE COVER           -7250.000 -7250.000 N DO 5 BY 1 STEP 40.000 0.000 ;
    CANNOTOCCUPY CORE            -5021.450 -4989.600 FS DO 100 BY 595 STEP 0.700 16.800 ;
    CANNOTOCCUPY CORE            -5021.450 -4998.000 N DO 100 BY 595 STEP 0.700 16.800 ;
    TRACKS X -6148.800 DO 17569 STEP 0.700 LAYER RX ;
    TRACKS Y -6148.800 DO 20497 STEP 0.600 LAYER RX ;

  FLOORPLAN 100%
    CANPLACE COVER           -7315.000 -7315.000 N DO 1 BY 1 STEP 0.000 0.000 ;
    CANPLACE COVER           -7250.000 -7250.000 N DO 5 BY 1 STEP 40.000 0.000 ;
    CANPLACE CORE            -5021.450 -4998.000 N DO 14346 BY 595 STEP 0.700 16.800 ;
    CANPLACE CORE            -5021.450 -4989.600 FS DO 14346 BY 595 STEP 0.700 16.800 ;
    CANNOTOCCUPY CORE            -5021.450 -4989.600 FS DO 100 BY 595 STEP 0.700 16.800 ;
    CANNOTOCCUPY CORE            -5021.450 -4998.000 N DO 100 BY 595 STEP 0.700 16.800 ;
  END 100%
  GCELLGRID X               -6157.200 DO 1467 STEP 8.400 ;
  GCELLGRID Y               -6157.200 DO 1467 STEP 8.400 ;
END M7E4XXX

MACRO CHK3A
	CLASS RING ;
        SOURCE USER ;
        FOREIGN CHKS 0 0 FN ;
        ORIGIN 0.9 0.9 ;
        EEQ CHK1 ; 
        LEQ CHK2 ; 
	SIZE 10.8 BY 28.8 ;
#  for testing the lefrWarning.log file
#        SITE CORE ;
	SYMMETRY X Y R90  ;
	SITE CORE ;
        POWER 1.0 ;
        PROPERTY stringProp "first" integerProp 1 WEIGHT 30.31 ;

	PIN GND
		TAPERRULE RULE1 ;
                FOREIGN GROUND ( 0 0 ) E ;
                LEQ  A ;
		DIRECTION INOUT ;
		USE GROUND ;
		SHAPE ABUTMENT ;
                INPUTNOISEMARGIN  6.1 2.3 ;
                OUTPUTNOISEMARGIN 5.0  4.6 ;
                OUTPUTRESISTANCE 7.4 5.4 ;
                POWER 2.0 ;
                LEAKAGE 1.0 ;
                CAPACITANCE 0.1 ;        
                RESISTANCE 0.2 ;
                PULLDOWNRES 0.5 ;
                TIEOFFR 0.8 ; 
                VHI 5 ;        
                VLO 0 ;        
                RISEVOLTAGETHRESHOLD 2.0 ;
                FALLVOLTAGETHRESHOLD 2.0 ;
                RISETHRESH 22 ;        
                FALLTHRESH 100 ;        
                RISESATCUR 4 ;        
                FALLSATCUR .5 ;        
                CURRENTSOURCE ACTIVE ;            
#               ANTENNASIZE 0.6 LAYER RX ;
#       	ANTENNAMETALAREA 3 LAYER M1 ;
#               ANTENNAMETALAREA 4 LAYER M2 ;
#               ANTENNAMETALLENGTH 5 LAYER M1 ;
#               ANTENNAMETALLENGTH 6 LAYER M2 ;
		RISESLEWLIMIT 0.01 ;
		FALLSLEWLIMIT 0.02 ;
                MAXDELAY 21 ;                        
		MAXLOAD 0.1 ;
		PROPERTY TYPE "special" intProp 23 realProp 24.25 ;
                IV_TABLES LOWT HIGHT ;

		PORT
                    CLASS CORE ;
	            LAYER M1 SPACING 0.05 ;
                         WIDTH 1.0 ;
			 RECT -0.9 3 9.9 6 ;
                    VIA 100 300 IN1X ;
		END
	END GND
	PIN VDD
		DIRECTION INOUT ;
                FOREIGN GROUND  STRUCTURE ( 0 0 ) E ;
		USE POWER ;
		SHAPE ABUTMENT ;
                PORT
                END
		PORT
                   CLASS NONE ;
		   LAYER M1 ;
			RECT ITERATE -0.9 21 9.9 24 
                            DO 1 BY 2 STEP 1 1 ;
                   VIA ITERATE 100 300 nd1VIA12 
                            DO 1 BY 2 STEP 1 2 ;
		END
#               ANTENNAMETALAREA 3 LAYER M1 ;
#               ANTENNAMETALAREA 4 LAYER M2 ;
#               ANTENNAMETALLENGTH 5 LAYER M1 ;
#               ANTENNAMETALLENGTH 6 LAYER M2 ;
                # Test for combination of both 5.3 & 5.4, which is not allowed
                # ANTENNAPARTIALMETALAREA 4 LAYER M1 ;
                LEAKAGE 1.0 ;
                FALLVOLTAGETHRESHOLD 2.0 ;
                RISEVOLTAGETHRESHOLD 2.0 ;
                CURRENTSOURCE ACTIVE ;
	END VDD
	PIN PA3
		DIRECTION INPUT ;
                # 5.4
                ANTENNAPARTIALMETALAREA 4 LAYER M1 ;
                ANTENNAPARTIALMETALAREA 5 LAYER M2 ;
                ANTENNAPARTIALMETALSIDEAREA 5 LAYER M2 ;
                ANTENNAPARTIALMETALSIDEAREA 6 LAYER M2 ;
                ANTENNAPARTIALMETALSIDEAREA 7 LAYER M2 ;
                ANTENNAGATEAREA 1 LAYER M1 ;
                ANTENNAGATEAREA 2 ;
                ANTENNAGATEAREA 3 LAYER M3 ;
                ANTENNADIFFAREA 1 LAYER M1 ;
                ANTENNAMAXAREACAR 1 LAYER L1 ;
                ANTENNAMAXAREACAR 2 LAYER L2 ;
                ANTENNAMAXAREACAR 3 LAYER L3 ;
                ANTENNAMAXAREACAR 4 LAYER L4 ;
                ANTENNAMAXSIDEAREACAR 1 LAYER L1 ;
                ANTENNAMAXSIDEAREACAR 2 LAYER L2 ;
                ANTENNAPARTIALCUTAREA 1 ;
                ANTENNAPARTIALCUTAREA 2 LAYER M2 ;
                ANTENNAPARTIALCUTAREA 3 ;
                ANTENNAPARTIALCUTAREA 4 LAYER M4 ;
                ANTENNAMAXCUTCAR 1 LAYER L1 ;
                ANTENNAMAXCUTCAR 2 LAYER L2 ;
                ANTENNAMAXCUTCAR 3 LAYER L3 ;
                # Test for combination of both 5.3 & 5.4, which is not allowed
		# ANTENNAMETALLENGTH 5 LAYER M1 ;
		PORT
			LAYER M1 SPACING 0.02 ;
			 RECT 1.35 -0.45 2.25 0.45 ;
			 RECT -0.45 -0.45 0.45 0.45 ;
		END
		PORT
			LAYER PC DESIGNRULEWIDTH 0.05 ;
			 RECT -0.45 12.15 0.45 13.05 ;
		END
		PORT
			LAYER PC ;
			 RECT -0.45 24.75 0.45 25.65 ;
		END
	END PA3
	PIN PA0
		DIRECTION INPUT ;
                MUSTJOIN PA3 ;
		PORT
                        CLASS NONE ;
			LAYER M1 ;
			 RECT 8.55 8.55 9.45 9.45 ;
			 RECT 6.75 6.75 7.65 7.65 ;
			 RECT 6.75 8.55 7.65 9.45 ;
			 RECT 6.75 10.35 7.65 11.25 ;
		END
		PORT
                        CLASS CORE ;
			LAYER PC ;
			 RECT 8.55 24.75 9.45 25.65 ;
		END
		PORT
			LAYER PC ;
			 RECT 6.75 1.35 7.65 2.25 ;
		END
		PORT
			LAYER PC ;
			 RECT 6.75 24.75 7.65 25.65 ;
		END
		PORT
			LAYER PC ;
			 RECT 4.95 1.35 5.85 2.25 ;
		END
	END PA0
	PIN PA1
		DIRECTION INPUT ;
		PORT
			LAYER M1 ;
			 RECT 8.55 -0.45 9.45 0.45 ;
			 RECT 6.75 -0.45 7.65 0.45 ;
		END
		PORT
			LAYER M1 ;
			 RECT 8.55 12.15 9.45 13.05 ;
			 RECT 6.75 12.15 7.65 13.05 ;
			 RECT 4.95 12.15 5.85 13.05 ;
		END
		PORT
			LAYER PC ;
			 RECT 4.95 24.75 5.85 25.65 ;
		END
		PORT
			LAYER PC ;
			 RECT 3.15 24.75 4.05 25.65 ;
		END
	END PA1
	PIN PA20
		DIRECTION INPUT ;
		PORT
			LAYER M1 ;
			 POLYGON 15 35 15 60 65 60 65 35 15 35 ;
		END
		PORT
			LAYER M1 ;
			 PATH 8.55 12.15 9.45 13.05 ;
		END
	END PA20
	PIN PA21
		DIRECTION OUTPUT TRISTATE ;
		PORT
			LAYER M1 ;
			POLYGON ITERATE 20 35 20 60 70 60 70 35
                                DO 1 BY 2 STEP 5 5 ;
		END
		PORT
			LAYER M1 ;
			PATH ITERATE 5.55 12.15 10.45 13.05 
                                 DO 1 BY 2 STEP 2 2 ;
		END
	END PA21
	OBS
		LAYER M1 SPACING 5.6 ;
		 RECT 6.6 -0.6 9.6 0.6 ;
		 RECT 4.8 12 9.6 13.2 ;
		 RECT 3 13.8 7.8 16.8 ;
		 RECT 3 -0.6 6 0.6 ;
		 RECT 3 8.4 6 11.4 ;
		 RECT 3 8.4 4.2 16.8 ;
		 RECT -0.6 13.8 4.2 16.8 ;
		 RECT -0.6 -0.6 2.4 0.6 ;
		 RECT 6.6 6.6 9.6 11.4 ;
		 RECT 6.6 6.6 7.8 11.4 ;
	END 
    TIMING
    FROMPIN PA21 ;
    TOPIN PA20 ;
    RISE INTRINSIC .39 .41 1.2 .25 .29 1.8 .67 .87 2.2
	 VARIABLE 0.12 0.13 ;
    FALL INTRINSIC .24 .29 1.3 .26 .31 1.7 .6 .8 2.1
	 VARIABLE 0.11 0.14 ;
    RISERS 83.178 90.109 ;
    FALLRS 76.246 97.041 ;
    RISECS 0.751 0.751 ;
    FALLCS 0.751 0.751 ;
    RISET0 0.65493 0.65493 ;
    FALLT0 0.38 0.38 ;
    RISESATT1 0 0 ;
    FALLSATT1 0.15 0.15 ;
    UNATENESS INVERT ;
   END TIMING
END CHK3A

MACRO INV

   CLASS CORE ;
   SOURCE BLOCK ;
   FOREIGN INVS ;
   POWER 1.0 ;
   SIZE 67.2 BY 24 ;
   SYMMETRY X Y R90 ;
   SITE CORE1 ;

   PIN Z DIRECTION OUTPUT ;
    USE SIGNAL ;
    RISETHRESH 22 ;
    FALLTHRESH 100 ;
    RISESATCUR 4 ;
    FALLSATCUR .5 ;
    VLO 0 ;
    VHI 5 ;
    CAPACITANCE 0.1 ;
    MAXDELAY 21 ;
    POWER 0.1 ;
    PORT
        LAYER M2 ;
           PATH 30.8 9 42 9 ;
    END
   END Z

   PIN A DIRECTION INPUT ;
    USE ANALOG ;
    RISETHRESH 22 ;
    FALLTHRESH 100 ;
    RISESATCUR 4 ;
    FALLSATCUR .5 ;
    VLO 0 ;
    VHI 5 ;
    CAPACITANCE 0.08 ;
    MAXDELAY 21 ;
    PORT
        LAYER M1 ;
           PATH 25.2 15 ;
    END
   END A

   PIN VDD DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    POWER 0.1 ;
    PORT
        LAYER M1 ;
           WIDTH 5.6 ;
           PATH 50.4 2.8 50.4 21.2 ;
    END
   END VDD

   PIN VSS DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    POWER 0.1 ;
    PORT
        LAYER M1 ;
           WIDTH 5.6 ;
           PATH 16.8 2.8 16.8 21.2 ;
    END
   END VSS

   TIMING
    FROMPIN A ;
    TOPIN Z ;
    RISE INTRINSIC .39 .41 1.2 .25 .29 1.8 .67 .87 2.2
         VARIABLE 0.12 0.13 ;
    FALL INTRINSIC .24 .29 1.3 .26 .31 1.7 .6 .8 2.1
         VARIABLE 0.11 0.14 ;
    RISERS 83.178 90.109 ;
    FALLRS 76.246 97.041 ;
    RISECS 0.751 0.751 ;
    FALLCS 0.751 0.751 ;
    RISET0 0.65493 0.65493 ;
    FALLT0 0.38 0.38 ;
    RISESATT1 0 0 ;
    FALLSATT1 0.15 0.15 ;
    UNATENESS INVERT ;
   END TIMING

   OBS
    LAYER M1 DESIGNRULEWIDTH 4.5 ;
        WIDTH 0.1 ;
        RECT 24.1 1.5 43.5 16.5 ;
        RECT ITERATE 24.1 1.5 43.5 16.5
             DO 2 BY 1 STEP 20.0 0 ;
        PATH ITERATE 532.0 534 1999.2 534
             DO 1 BY 2 STEP 0 1446 ;
        VIA ITERATE 470.4 475 VIABIGPOWER12
             DO 2 BY 2 STEP 1590.4 1565 ;
        PATH 532.0 534 1999.2 534 ;
        PATH 532.0 1980 1999.2 1980 ;
        VIA 470.4 475 VIABIGPOWER12 ;
        VIA 2060.8 475 VIABIGPOWER12 ;
        VIA 470.4 2040 VIABIGPOWER12 ;
        VIA 2060.8 2040 VIABIGPOWER12 ;
        RECT 44.1 1.5 63.5 16.5 ;
   END

END INV

MACRO INV_B
   EEQ INV ;

   CLASS CORE SPACER ;
   FOREIGN INVS ( 4 5 ) ;
   POWER 1.0 ;
   SIZE 67.2 BY 24 ;
   SYMMETRY X Y R90 ;
   SITE CORE1 ;
   PIN Z DIRECTION OUTPUT ;
    USE CLOCK ;
    RISETHRESH 22 ;
    FALLTHRESH 100 ;
    RISESATCUR 4 ;
    FALLSATCUR .5 ;
    VLO 0 ;
    VHI 5 ;
    CAPACITANCE 0.1 ;
    MAXDELAY 21 ;
    POWER 0.1 ;
    PORT
        LAYER M2 ;
           PATH 30.8 9 42 9 ;
    END
   END Z

   PIN A DIRECTION FEEDTHRU ;
    USE SIGNAL ;
    RISETHRESH 22 ;
    FALLTHRESH 100 ;
    RISESATCUR 4 ;
    FALLSATCUR .5 ;
    VLO 0 ;
    VHI 5 ;
    CAPACITANCE 0.08 ;
    MAXDELAY 21 ;
    PORT
        LAYER M1 ;
           PATH 25.2 15 ;
    END
   END A

   PIN VDD DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    POWER 0.1 ;
    PORT
        LAYER M1 ;
           WIDTH 5.6 ;
           PATH 50.4 2.8 50.4 21.2 ;
    END
   END VDD

   PIN VSS DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    POWER 0.1 ;
    PORT
        LAYER M1 ;
           WIDTH 5.6 ;
           PATH 16.8 2.8 16.8 21.2 ;
    END
   END VSS

   TIMING
    FROMPIN A ;
    TOPIN Z ;
    RISE INTRINSIC .39 .41 1.2 .25 .29 1.8 .67 .87 2.2
        VARIABLE 0.12 0.13 ;
    FALL INTRINSIC .24 .29 1.3 .26 .31 1.7 .6 .8 2.1
        VARIABLE 0.11 0.14 ;
    RISERS 83.178 90.109 ;
    FALLRS 76.246 97.041 ;
    RISECS 0.751 0.751 ;
    FALLCS 0.751 0.751 ;
    RISET0 0.65493 0.65493 ;
    FALLT0 0.38 0.38 ;
    RISESATT1 0 0 ;
    FALLSATT1 0.15 0.15 ;
    UNATENESS INVERT ;
   END TIMING

   OBS
    LAYER M1 ;
        RECT 24.1 1.5 43.5 16.5 ;
   END

END INV_B

MACRO DFF3

   CLASS CORE ANTENNACELL ;
   FOREIGN DFF3S ;
   POWER 4.0 ;
   SIZE 67.2 BY 210 ;
   SYMMETRY X Y R90 ;
   SITE CORE 34 54 FE DO 30 BY 3 STEP 1 1 ;
   SITE CORE1 21 68 S DO 30 BY 3 STEP 2 2 ;

   PIN Q DIRECTION OUTPUT ;
    USE SIGNAL ;
    RISETHRESH 22 ;
    FALLTHRESH 100 ;
    RISESATCUR 4 ;
    FALLSATCUR .5 ;
    VLO 0 ;
    VHI 5 ;
    CAPACITANCE 0.12 ;
    MAXDELAY 20 ;
    POWER 0.4 ;
    PORT
        LAYER M2 ;
           PATH 19.6 99 47.6 99 ;
    END
   END Q

   PIN QN DIRECTION OUTPUT ;
    USE SIGNAL ;
    RISETHRESH 22 ;
    FALLTHRESH 100 ;
    RISESATCUR 4 ;
    FALLSATCUR .5 ;
    VLO 0 ;
    VHI 5 ;
    CAPACITANCE 0.11 ;
    MAXDELAY 20 ;
    POWER 0.4 ;
    PORT
        LAYER M2 ;
           PATH 25.2 123 42 123 ;
    END
   END QN

   PIN D DIRECTION INPUT ;
    USE SIGNAL ;
    RISETHRESH 22 ;
    FALLTHRESH 100 ;
    RISESATCUR 4 ;
    FALLSATCUR .5 ;
    VLO 0 ;
    VHI 5 ;
    CAPACITANCE 0.13 ;
    MAXDELAY 20 ;
    POWER 0.4 ;
    PORT
        LAYER M1 ;
           PATH 30.8 51 ;
    END
   END D

   PIN G DIRECTION INPUT ;
    USE SIGNAL ;
    RISETHRESH 22 ;
    FALLTHRESH 100 ;
    RISESATCUR 4 ;
    FALLSATCUR .5 ;
    VLO 0 ;
    VHI 5 ;
    CAPACITANCE 0.11 ;
    MAXDELAY 20 ;
    POWER 0.4 ;
    PORT
        LAYER M1 ;
           PATH 25.2 3 ;
    END
   END G

   PIN CD DIRECTION INPUT ;
    USE CLOCK ;
    RISETHRESH 22 ;
    FALLTHRESH 100 ;
    RISESATCUR 4 ;
    FALLSATCUR .5 ;
    VLO 0 ;
    VHI 5 ;
    CAPACITANCE 0.1 ;
    MAXDELAY 20 ;
    POWER 0.4 ;
    PORT
        LAYER M1 ;
           PATH 36.4 75 ;
    END
   END CD

   PIN VDD DIRECTION INOUT ;
    SHAPE RING ;
    POWER 0.4 ;
    PORT
        LAYER M1 ;
           WIDTH 5.6 ;
           PATH 50.4 2.8 50.4 207.2 ;
    END
   END VDD

   PIN VSS DIRECTION INOUT ;
    SHAPE FEEDTHRU ;
    POWER 0.4 ;
    PORT
        LAYER M1 ;
           WIDTH 5.6 ;
           PATH 16.8 2.8 16.8 207.2 ;
    END
   END VSS

   TIMING
    FROMPIN D ;
    TOPIN Q ;
    RISE INTRINSIC .51 .6 1.4 .37 .45 1.7 .6 .81 2.1
        VARIABLE 0.06 0.1 ;
    FALL INTRINSIC 1 1.2 1.4 1.77 1.85 1.8 .56 .81 2.4
        VARIABLE 0.08 0.09 ;
    RISERS 41.589 69.315 ;
    FALLRS 55.452 62.383 ;
    RISECS 0.113 0.113 ;
    FallCS 0.113 0.113 ;
    RISET0 0.023929 0.023929 ;
    FALLT0 0.38 0.38 ;
    RISESATT1 0 0 ;
    FALLSATT1 0.15 0.15 ;
    UNATENESS      NONINVERT ;
   END TIMING

   OBS
    LAYER M1 DESIGNRULEWIDTH 0.15 ;
        RECT 24.1 1.5 43.5 208.5 ;
        PATH 8.4 3 8.4 123 ;
        PATH 58.8 3 58.8 123 ;
        PATH 64.4 3 64.4 123 ;
   END

END DFF3

MACRO BUF1
  CLASS ENDCAP BOTTOMLEFT ;
  PIN IN
    ANTENNAGATEAREA 1 ;
    ANTENNAGATEAREA 3 ;
    ANTENNADIFFAREA 0 ;
    ANTENNAMODEL OXIDE2 ;
    ANTENNAGATEAREA 2 ;
    ANTENNAGATEAREA 4 ;
    ANTENNADIFFAREA 0 ;
  END IN
  PIN IN2
    ANTENNAGATEAREA 1 ;
  END IN2
  PIN IN3
    SHAPE ABUTMENT ;
  END IN3
END BUF1

MACRO DFF4
   CLASS COVER BUMP ;
   FOREIGN DFF3S ;
   POWER 4.0 ;
END DFF4

MACRO DFF5
   CLASS COVER ;
   FOREIGN DFF3S ;
END DFF5

MACRO mydriver
   CLASS PAD AREAIO ;
   FOREIGN DFF3S ;
END mydriver

MACRO myblackbox
   CLASS BLOCK BLACKBOX ;
   FOREIGN DFF3S ;
END myblackbox

ANTENNAINPUTGATEAREA 45 ;
ANTENNAINOUTDIFFAREA 65 ;
ANTENNAOUTPUTDIFFAREA 55 ;

#INPUTPINANTENNASIZE 1 ;
#OUTPUTPINANTENNASIZE -1 ;
#INOUTPINANTENNASIZE -1 ;

BEGINEXT "SIGNATURE"
	CREATOR "CADENCE"
	DATE "04/14/98"
ENDEXT

END LIBRARY
